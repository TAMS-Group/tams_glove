// 2023-2024 Philipp Ruppel

`include "tac_baseline.sv"
`include "tac_test_inc.sv"