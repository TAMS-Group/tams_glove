// 2023-2024 Philipp Ruppel

`include "tac_new.v"
`include "tac_test_inc.sv"