// 2023-2024 Philipp Ruppel

`include "shfloat.v"
