// 2023-2024 Philipp Ruppel

`include "tac_old.v"
`include "tac_test_inc.sv"